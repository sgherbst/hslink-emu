`timescale 1ns/1ps

package globals;

    parameter ROM_DIR_PATH = "/horowitz/users/sherbst/msemu/build/roms/";

endpackage // globals
