package iotype;

	typedef real voltage_t;

endpackage
