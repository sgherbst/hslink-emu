`timescale 1ns/1ps

package globals;

    parameter ROM_DIR_PATH = "//Mac/Home/Desktop/msemu/build/roms/";

endpackage // globals
