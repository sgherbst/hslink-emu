module buff import iotype::*; (
	input voltage_t x,
	output voltage_t y
); 

	assign y = x;

endmodule
